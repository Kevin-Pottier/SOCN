
Library IEEE;
 use IEEE.std_logic_1164.all;

package PkgS51Timer is

 type T_TIMERSM is (TM_IDLE, TM_DECR, TM_RELOAD);

end PkgS51Timer;

package body PkgS51Timer is

end;

