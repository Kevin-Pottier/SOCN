
----------------------------------------------------------------
-- 
-- DATE CREATED :    Tue Aug  6 2006
-- 
-- LIBRARY      :    c35_CORELIB_3B
-- REVISION     :    2.1 bka
-- TECHNOLOGY   :    cmos
-- TIME SCALE   :    1 ps
-- LOGIC SYSTEM :    IEEE-1164
-- NOTES        :    VITAL, TimingChecksOn(TRUE), XGenerationOn(TRUE), TimingMessage(TRUE), OnEvent 
--                   Owner: austriamicrosystems AG  HIT-Kit: Digital
-- HISTORY      :
-- 
----------------------------------------------------------------

----- CELL ADD21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ADD21_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ADD21_3B : entity is TRUE;
end ADD21_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of ADD21_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (A_ipd) AND (B_ipd);
      S_zd := (A_ipd) XOR (B_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_ADD21_VITAL of ADD21_3B is
   for VITAL
   end for;
end CFG_ADD21_VITAL;


----- CELL ADD22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ADD22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ADD22_3B : entity is TRUE;
end ADD22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of ADD22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (A_ipd) AND (B_ipd);
      S_zd := (A_ipd) XOR (B_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_ADD22_VITAL of ADD22_3B is
   for VITAL
   end for;
end CFG_ADD22_VITAL;


----- CELL ADD31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ADD31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_CI_CO                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_CI_S                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_CI                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ADD31_3B : entity is TRUE;
end ADD31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of ADD31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd :=
       ((A_ipd) AND (CI_ipd)) OR ((B_ipd) AND (CI_ipd)) OR ((A_ipd) AND
         (B_ipd));
      S_zd := (B_ipd) XOR (CI_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (CI_ipd'last_event, tpd_CI_CO, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (CI_ipd'last_event, tpd_CI_S, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_ADD31_VITAL of ADD31_3B is
   for VITAL
   end for;
end CFG_ADD31_VITAL;


----- CELL ADD32 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ADD32_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_CO                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_CI_CO                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_S                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_CI_S                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_CI                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ADD32_3B : entity is TRUE;
end ADD32_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of ADD32_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd :=
       ((A_ipd) AND (CI_ipd)) OR ((B_ipd) AND (CI_ipd)) OR ((A_ipd) AND
         (B_ipd));
      S_zd := (B_ipd) XOR (CI_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (CI_ipd'last_event, tpd_CI_CO, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (CI_ipd'last_event, tpd_CI_S, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_ADD32_VITAL of ADD32_3B is
   for VITAL
   end for;
end CFG_ADD32_VITAL;


----- CELL AOI210 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI210_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI210_3B : entity is TRUE;
end AOI210_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI210_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI210_VITAL of AOI210_3B is
   for VITAL
   end for;
end CFG_AOI210_VITAL;


----- CELL AOI211 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI211_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI211_3B : entity is TRUE;
end AOI211_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI211_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI211_VITAL of AOI211_3B is
   for VITAL
   end for;
end CFG_AOI211_VITAL;


----- CELL AOI212 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI212_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI212_3B : entity is TRUE;
end AOI212_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI212_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI212_VITAL of AOI212_3B is
   for VITAL
   end for;
end CFG_AOI212_VITAL;


----- CELL AOI220 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI220_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI220_3B : entity is TRUE;
end AOI220_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI220_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((C_ipd) AND (D_ipd)) OR ((A_ipd) AND (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI220_VITAL of AOI220_3B is
   for VITAL
   end for;
end CFG_AOI220_VITAL;


----- CELL AOI221 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI221_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI221_3B : entity is TRUE;
end AOI221_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI221_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((C_ipd) AND (D_ipd)) OR ((A_ipd) AND (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI221_VITAL of AOI221_3B is
   for VITAL
   end for;
end CFG_AOI221_VITAL;


----- CELL AOI222 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI222_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI222_3B : entity is TRUE;
end AOI222_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI222_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((C_ipd) AND (D_ipd)) OR ((A_ipd) AND (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI222_VITAL of AOI222_3B is
   for VITAL
   end for;
end CFG_AOI222_VITAL;


----- CELL AOI310 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI310_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI310_3B : entity is TRUE;
end AOI310_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI310_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((D_ipd) OR ((A_ipd) AND (B_ipd) AND (C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI310_VITAL of AOI310_3B is
   for VITAL
   end for;
end CFG_AOI310_VITAL;


----- CELL AOI311 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI311_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI311_3B : entity is TRUE;
end AOI311_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI311_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((D_ipd) OR ((A_ipd) AND (B_ipd) AND (C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI311_VITAL of AOI311_3B is
   for VITAL
   end for;
end CFG_AOI311_VITAL;


----- CELL AOI312 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI312_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI312_3B : entity is TRUE;
end AOI312_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI312_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((D_ipd) OR ((A_ipd) AND (B_ipd) AND (C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI312_VITAL of AOI312_3B is
   for VITAL
   end for;
end CFG_AOI312_VITAL;


----- CELL AOI2110 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI2110_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI2110_3B : entity is TRUE;
end AOI2110_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI2110_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR (D_ipd) OR ((A_ipd) AND (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI2110_VITAL of AOI2110_3B is
   for VITAL
   end for;
end CFG_AOI2110_VITAL;


----- CELL AOI2111 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI2111_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI2111_3B : entity is TRUE;
end AOI2111_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI2111_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR (D_ipd) OR ((A_ipd) AND (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI2111_VITAL of AOI2111_3B is
   for VITAL
   end for;
end CFG_AOI2111_VITAL;


----- CELL AOI2112 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI2112_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI2112_3B : entity is TRUE;
end AOI2112_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of AOI2112_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR (D_ipd) OR ((A_ipd) AND (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_AOI2112_VITAL of AOI2112_3B is
   for VITAL
   end for;
end CFG_AOI2112_VITAL;


----- CELL BUF2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUF2_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUF2_3B : entity is TRUE;
end BUF2_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUF2_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_BUF2_VITAL of BUF2_3B is
   for VITAL
   end for;
end CFG_BUF2_VITAL;


----- CELL BUF4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUF4_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUF4_3B : entity is TRUE;
end BUF4_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUF4_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_BUF4_VITAL of BUF4_3B is
   for VITAL
   end for;
end CFG_BUF4_VITAL;


----- CELL BUF6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUF6_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUF6_3B : entity is TRUE;
end BUF6_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUF6_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_BUF6_VITAL of BUF6_3B is
   for VITAL
   end for;
end CFG_BUF6_VITAL;


----- CELL BUF8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUF8_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUF8_3B : entity is TRUE;
end BUF8_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUF8_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_BUF8_VITAL of BUF8_3B is
   for VITAL
   end for;
end CFG_BUF8_VITAL;


----- CELL BUF12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUF12_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUF12_3B : entity is TRUE;
end BUF12_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUF12_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_BUF12_VITAL of BUF12_3B is
   for VITAL
   end for;
end CFG_BUF12_VITAL;


----- CELL BUF15 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUF15_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUF15_3B : entity is TRUE;
end BUF15_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUF15_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_BUF15_VITAL of BUF15_3B is
   for VITAL
   end for;
end CFG_BUF15_VITAL;


----- CELL BUFE2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFE2_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_E_Q                        :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFE2_3B : entity is TRUE;
end BUFE2_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFE2_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFE2_VITAL of BUFE2_3B is
   for VITAL
   end for;
end CFG_BUFE2_VITAL;


----- CELL BUFE4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFE4_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_E_Q                        :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFE4_3B : entity is TRUE;
end BUFE4_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFE4_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFE4_VITAL of BUFE4_3B is
   for VITAL
   end for;
end CFG_BUFE4_VITAL;


----- CELL BUFE6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFE6_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_E_Q                        :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFE6_3B : entity is TRUE;
end BUFE6_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFE6_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFE6_VITAL of BUFE6_3B is
   for VITAL
   end for;
end CFG_BUFE6_VITAL;


----- CELL BUFE8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFE8_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_E_Q                        :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFE8_3B : entity is TRUE;
end BUFE8_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFE8_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFE8_VITAL of BUFE8_3B is
   for VITAL
   end for;
end CFG_BUFE8_VITAL;


----- CELL BUFE10 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFE10_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_E_Q                        :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFE10_3B : entity is TRUE;
end BUFE10_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFE10_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFE10_VITAL of BUFE10_3B is
   for VITAL
   end for;
end CFG_BUFE10_VITAL;


----- CELL BUFE12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFE12_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_E_Q                        :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFE12_3B : entity is TRUE;
end BUFE12_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFE12_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFE12_VITAL of BUFE12_3B is
   for VITAL
   end for;
end CFG_BUFE12_VITAL;


----- CELL BUFE15 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFE15_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_E_Q                        :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFE15_3B : entity is TRUE;
end BUFE15_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFE15_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (E_ipd'last_event, VitalExtendToFillDelay(tpd_E_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFE15_VITAL of BUFE15_3B is
   for VITAL
   end for;
end CFG_BUFE15_VITAL;


----- CELL BUFT2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFT2_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_EN_Q                       :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_EN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      EN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFT2_3B : entity is TRUE;
end BUFT2_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFT2_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, EN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (EN_ipd'last_event, VitalExtendToFillDelay(tpd_EN_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFT2_VITAL of BUFT2_3B is
   for VITAL
   end for;
end CFG_BUFT2_VITAL;


----- CELL BUFT4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFT4_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_EN_Q                       :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_EN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      EN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFT4_3B : entity is TRUE;
end BUFT4_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFT4_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, EN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (EN_ipd'last_event, VitalExtendToFillDelay(tpd_EN_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFT4_VITAL of BUFT4_3B is
   for VITAL
   end for;
end CFG_BUFT4_VITAL;


----- CELL BUFT6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFT6_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_EN_Q                       :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_EN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      EN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFT6_3B : entity is TRUE;
end BUFT6_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFT6_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, EN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (EN_ipd'last_event, VitalExtendToFillDelay(tpd_EN_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFT6_VITAL of BUFT6_3B is
   for VITAL
   end for;
end CFG_BUFT6_VITAL;


----- CELL BUFT8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFT8_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_EN_Q                       :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_EN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      EN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFT8_3B : entity is TRUE;
end BUFT8_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFT8_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, EN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (EN_ipd'last_event, VitalExtendToFillDelay(tpd_EN_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFT8_VITAL of BUFT8_3B is
   for VITAL
   end for;
end CFG_BUFT8_VITAL;


----- CELL BUFT10 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFT10_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_EN_Q                       :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_EN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      EN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFT10_3B : entity is TRUE;
end BUFT10_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFT10_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, EN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (EN_ipd'last_event, VitalExtendToFillDelay(tpd_EN_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFT10_VITAL of BUFT10_3B is
   for VITAL
   end for;
end CFG_BUFT10_VITAL;


----- CELL BUFT12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFT12_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_EN_Q                       :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_EN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      EN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFT12_3B : entity is TRUE;
end BUFT12_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFT12_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, EN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (EN_ipd'last_event, VitalExtendToFillDelay(tpd_EN_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFT12_VITAL of BUFT12_3B is
   for VITAL
   end for;
end CFG_BUFT12_VITAL;


----- CELL BUFT15 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFT15_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_EN_Q                       :	VitalDelayType01z := 
               (1 ps, 1 ps, 1 ps, 1 ps, 1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_EN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      EN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFT15_3B : entity is TRUE;
end BUFT15_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUFT15_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL EN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (EN_ipd, EN, tipd_EN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, EN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalBUFIF0 (data => A_ipd,
              enable => EN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, VitalExtendToFillDelay(tpd_A_Q), TRUE),
                 1 => (EN_ipd'last_event, VitalExtendToFillDelay(tpd_EN_Q), TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL;

configuration CFG_BUFT15_VITAL of BUFT15_3B is
   for VITAL
   end for;
end CFG_BUFT15_VITAL;


----- CELL BUSHD -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUSHD_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	inout STD_ULOGIC := 'Z');
attribute VITAL_LEVEL0 of BUSHD_3B : entity is TRUE;
end BUSHD_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of BUSHD_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A)


   -- functionality results
   VARIABLE A_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE A_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
   A_zd := VitalBUF ( A, ('W', 'W', 'L', 'H'));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => A,
       GlitchData => A_GlitchData,
       OutSignalName => "A",
       OutTemp => A_zd,
       Paths => (0=>(A'last_event, VitalZeroDelay01Z, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);


end process;

end VITAL;

configuration CFG_BUSHD_VITAL of BUSHD_3B is
   for VITAL
   end for;
end CFG_BUSHD_VITAL;


----- CELL CLKBU2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBU2_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBU2_3B : entity is TRUE;
end CLKBU2_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKBU2_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKBU2_VITAL of CLKBU2_3B is
   for VITAL
   end for;
end CFG_CLKBU2_VITAL;


----- CELL CLKBU4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBU4_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBU4_3B : entity is TRUE;
end CLKBU4_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKBU4_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKBU4_VITAL of CLKBU4_3B is
   for VITAL
   end for;
end CFG_CLKBU4_VITAL;


----- CELL CLKBU6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBU6_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBU6_3B : entity is TRUE;
end CLKBU6_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKBU6_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKBU6_VITAL of CLKBU6_3B is
   for VITAL
   end for;
end CFG_CLKBU6_VITAL;


----- CELL CLKBU8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBU8_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBU8_3B : entity is TRUE;
end CLKBU8_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKBU8_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKBU8_VITAL of CLKBU8_3B is
   for VITAL
   end for;
end CFG_CLKBU8_VITAL;


----- CELL CLKBU12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBU12_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBU12_3B : entity is TRUE;
end CLKBU12_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKBU12_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKBU12_VITAL of CLKBU12_3B is
   for VITAL
   end for;
end CFG_CLKBU12_VITAL;


----- CELL CLKBU15 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBU15_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBU15_3B : entity is TRUE;
end CLKBU15_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKBU15_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKBU15_VITAL of CLKBU15_3B is
   for VITAL
   end for;
end CFG_CLKBU15_VITAL;


----- CELL CLKIN0 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN0_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN0_3B : entity is TRUE;
end CLKIN0_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN0_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN0_VITAL of CLKIN0_3B is
   for VITAL
   end for;
end CFG_CLKIN0_VITAL;


----- CELL CLKIN1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN1_3B : entity is TRUE;
end CLKIN1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN1_VITAL of CLKIN1_3B is
   for VITAL
   end for;
end CFG_CLKIN1_VITAL;


----- CELL CLKIN2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN2_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN2_3B : entity is TRUE;
end CLKIN2_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN2_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN2_VITAL of CLKIN2_3B is
   for VITAL
   end for;
end CFG_CLKIN2_VITAL;


----- CELL CLKIN3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN3_3B : entity is TRUE;
end CLKIN3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN3_VITAL of CLKIN3_3B is
   for VITAL
   end for;
end CFG_CLKIN3_VITAL;


----- CELL CLKIN4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN4_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN4_3B : entity is TRUE;
end CLKIN4_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN4_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN4_VITAL of CLKIN4_3B is
   for VITAL
   end for;
end CFG_CLKIN4_VITAL;


----- CELL CLKIN6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN6_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN6_3B : entity is TRUE;
end CLKIN6_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN6_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN6_VITAL of CLKIN6_3B is
   for VITAL
   end for;
end CFG_CLKIN6_VITAL;


----- CELL CLKIN8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN8_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN8_3B : entity is TRUE;
end CLKIN8_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN8_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN8_VITAL of CLKIN8_3B is
   for VITAL
   end for;
end CFG_CLKIN8_VITAL;


----- CELL CLKIN10 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN10_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN10_3B : entity is TRUE;
end CLKIN10_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN10_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN10_VITAL of CLKIN10_3B is
   for VITAL
   end for;
end CFG_CLKIN10_VITAL;


----- CELL CLKIN12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN12_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN12_3B : entity is TRUE;
end CLKIN12_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN12_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN12_VITAL of CLKIN12_3B is
   for VITAL
   end for;
end CFG_CLKIN12_VITAL;


----- CELL CLKIN15 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKIN15_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKIN15_3B : entity is TRUE;
end CLKIN15_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of CLKIN15_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_CLKIN15_VITAL of CLKIN15_3B is
   for VITAL
   end for;
end CFG_CLKIN15_VITAL;


----- CELL DF1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1_3B : entity is TRUE;
end DF1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DF1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               C_delayed, D_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DF1_VITAL of DF1_3B is
   for VITAL
   end for;
end CFG_DF1_VITAL;


----- CELL DF3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF3_3B : entity is TRUE;
end DF3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DF3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               C_delayed, D_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DF3_VITAL of DF3_3B is
   for VITAL
   end for;
end CFG_DF3_VITAL;


----- CELL DFC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1_3B : entity is TRUE;
end DFC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, D_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFC1_VITAL of DFC1_3B is
   for VITAL
   end for;
end CFG_DFC1_VITAL;


----- CELL DFC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC3_3B : entity is TRUE;
end DFC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, D_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFC3_VITAL of DFC3_3B is
   for VITAL
   end for;
end CFG_DFC3_VITAL;


----- CELL DFCP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFCP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFCP1_3B : entity is TRUE;
end DFCP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFCP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, D_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, RN_ipd, D_delayed, C_ipd));
      QN_zd := Violation XOR QN_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFCP1_VITAL of DFCP1_3B is
   for VITAL
   end for;
end CFG_DFCP1_VITAL;


----- CELL DFCP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFCP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFCP3_3B : entity is TRUE;
end DFCP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFCP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, D_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, RN_ipd, D_delayed, C_ipd));
      QN_zd := Violation XOR QN_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFCP3_VITAL of DFCP3_3B is
   for VITAL
   end for;
end CFG_DFCP3_VITAL;


----- CELL DFE1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1_3B : entity is TRUE;
end DFE1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFE1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1_Q_tab,
        DataIn => (
               C_delayed, Q_zd, D_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFE1_VITAL of DFE1_3B is
   for VITAL
   end for;
end CFG_DFE1_VITAL;


----- CELL DFE3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3_3B : entity is TRUE;
end DFE3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFE3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1_Q_tab,
        DataIn => (
               C_delayed, Q_zd, D_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFE3_VITAL of DFE3_3B is
   for VITAL
   end for;
end CFG_DFE3_VITAL;


----- CELL DFEC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEC1_3B : entity is TRUE;
end DFEC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFEC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, Q_zd, D_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFEC1_VITAL of DFEC1_3B is
   for VITAL
   end for;
end CFG_DFEC1_VITAL;


----- CELL DFEC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEC3_3B : entity is TRUE;
end DFEC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFEC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, Q_zd, D_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFEC3_VITAL of DFEC3_3B is
   for VITAL
   end for;
end CFG_DFEC3_VITAL;


----- CELL DFECP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFECP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFECP1_3B : entity is TRUE;
end DFECP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFECP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, E_delayed, Q_zd, D_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, Q_zd, D_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFECP1_VITAL of DFECP1_3B is
   for VITAL
   end for;
end CFG_DFECP1_VITAL;


----- CELL DFECP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFECP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFECP3_3B : entity is TRUE;
end DFECP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFECP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, E_delayed, Q_zd, D_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, Q_zd, D_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFECP3_VITAL of DFECP3_3B is
   for VITAL
   end for;
end CFG_DFECP3_VITAL;


----- CELL DFEP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEP1_3B : entity is TRUE;
end DFEP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFEP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFEP1_Q_tab,
        DataIn => (
               C_delayed, Q_zd, D_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFEP1_VITAL of DFEP1_3B is
   for VITAL
   end for;
end CFG_DFEP1_VITAL;


----- CELL DFEP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEP3_3B : entity is TRUE;
end DFEP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFEP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFEP1_Q_tab,
        DataIn => (
               C_delayed, Q_zd, D_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFEP3_VITAL of DFEP3_3B is
   for VITAL
   end for;
end CFG_DFEP3_VITAL;


----- CELL DFP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1_3B : entity is TRUE;
end DFP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               C_delayed, D_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFP1_VITAL of DFP1_3B is
   for VITAL
   end for;
end CFG_DFP1_VITAL;


----- CELL DFP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := -1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP3_3B : entity is TRUE;
end DFP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               C_delayed, D_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFP3_VITAL of DFP3_3B is
   for VITAL
   end for;
end CFG_DFP3_VITAL;


----- CELL DFS1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFS1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFS1_3B : entity is TRUE;
end DFS1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFS1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => 0 ps,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => 0 ps,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFS1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, D_delayed, SE_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFS1_VITAL of DFS1_3B is
   for VITAL
   end for;
end CFG_DFS1_VITAL;


----- CELL DFS3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFS3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFS3_3B : entity is TRUE;
end DFS3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFS3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFS1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, D_delayed, SE_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFS3_VITAL of DFS3_3B is
   for VITAL
   end for;
end CFG_DFS3_VITAL;


----- CELL DFSC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSC1_3B : entity is TRUE;
end DFSC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, D_delayed, SE_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSC1_VITAL of DFSC1_3B is
   for VITAL
   end for;
end CFG_DFSC1_VITAL;


----- CELL DFSC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSC3_3B : entity is TRUE;
end DFSC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, D_delayed, SE_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSC3_VITAL of DFSC3_3B is
   for VITAL
   end for;
end CFG_DFSC3_VITAL;


----- CELL DFSCP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSCP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSCP1_3B : entity is TRUE;
end DFSCP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSCP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, D_delayed, SE_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFSCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, SE_delayed, SD_delayed, D_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSCP1_VITAL of DFSCP1_3B is
   for VITAL
   end for;
end CFG_DFSCP1_VITAL;


----- CELL DFSCP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSCP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSCP3_3B : entity is TRUE;
end DFSCP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSCP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, D_delayed, SE_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFSCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, SE_delayed, SD_delayed, D_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSCP3_VITAL of DFSCP3_3B is
   for VITAL
   end for;
end CFG_DFSCP3_VITAL;


----- CELL DFSE1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSE1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSE1_3B : entity is TRUE;
end DFSE1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSE1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSE1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSE1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSE1_VITAL of DFSE1_3B is
   for VITAL
   end for;
end CFG_DFSE1_VITAL;


----- CELL DFSE3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSE3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSE3_3B : entity is TRUE;
end DFSE3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSE3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSE3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSE1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSE3_VITAL of DFSE3_3B is
   for VITAL
   end for;
end CFG_DFSE3_VITAL;


----- CELL DFSEC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSEC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSEC1_3B : entity is TRUE;
end DFSEC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSEC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSEC1_VITAL of DFSEC1_3B is
   for VITAL
   end for;
end CFG_DFSEC1_VITAL;


----- CELL DFSEC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSEC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 0 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSEC3_3B : entity is TRUE;
end DFSEC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSEC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSEC3_VITAL of DFSEC3_3B is
   for VITAL
   end for;
end CFG_DFSEC3_VITAL;


----- CELL DFSECP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSECP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSECP1_3B : entity is TRUE;
end DFSECP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSECP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFSECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, SE_delayed, E_delayed, Q_zd, D_delayed, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSECP1_VITAL of DFSECP1_3B is
   for VITAL
   end for;
end CFG_DFSECP1_VITAL;


----- CELL DFSECP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSECP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSECP3_3B : entity is TRUE;
end DFSECP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSECP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Tviol_RN_C_posedge or Pviol_C or Pviol_RN or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFSECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, SE_delayed, E_delayed, Q_zd, D_delayed, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSECP3_VITAL of DFSECP3_3B is
   for VITAL
   end for;
end CFG_DFSECP3_VITAL;


----- CELL DFSEP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSEP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSEP1_3B : entity is TRUE;
end DFSEP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSEP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSEP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSEP1_VITAL of DFSEP1_3B is
   for VITAL
   end for;
end CFG_DFSEP1_VITAL;


----- CELL DFSEP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSEP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_E_C_posedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSEP3_3B : entity is TRUE;
end DFSEP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSEP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, E_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Tviol_E_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSEP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, Q_zd, D_delayed, SE_delayed, E_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSEP3_VITAL of DFSEP3_3B is
   for VITAL
   end for;
end CFG_DFSEP3_VITAL;


----- CELL DFSP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSP1_3B : entity is TRUE;
end DFSP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, D_delayed, SE_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSP1_VITAL of DFSP1_3B is
   for VITAL
   end for;
end CFG_DFSP1_VITAL;


----- CELL DFSP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFSP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_D_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_D_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_D_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DFSP3_3B : entity is TRUE;
end DFSP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DFSP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, D_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_C_posedge,
          TimingData              => Tmkr_D_C_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_C_posedge_posedge,
          SetupLow                => tsetup_D_C_negedge_posedge,
          HoldHigh                => thold_D_C_posedge_posedge,
          HoldLow                 => thold_D_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_C_posedge or Pviol_C or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFSP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, D_delayed, SE_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      D_delayed := D_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DFSP3_VITAL of DFSP3_3B is
   for VITAL
   end for;
end CFG_DFSP3_VITAL;


----- CELL DL1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1_3B : entity is TRUE;
end DL1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DL1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Pviol_GN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DL1_VITAL of DL1_3B is
   for VITAL
   end for;
end CFG_DL1_VITAL;


----- CELL DL3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL3_3B : entity is TRUE;
end DL3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DL3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Pviol_GN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DL3_VITAL of DL3_3B is
   for VITAL
   end for;
end CFG_DL3_VITAL;


----- CELL DLC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := -1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1_3B : entity is TRUE;
end DLC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Pviol_GN or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLC1_VITAL of DLC1_3B is
   for VITAL
   end for;
end CFG_DLC1_VITAL;


----- CELL DLC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := -1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC3_3B : entity is TRUE;
end DLC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Pviol_GN or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLC3_VITAL of DLC3_3B is
   for VITAL
   end for;
end CFG_DLC3_VITAL;


----- CELL DLCP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := -1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := -1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCP1_3B : entity is TRUE;
end DLCP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLCP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DLCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Tviol_SN_GN_posedge or Pviol_RN or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLCP1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLCP1_QN_tab,
        DataIn => (
               SN_ipd, GN_ipd, RN_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 3 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 3 => (SN_ipd'last_event, tpd_SN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLCP1_VITAL of DLCP1_3B is
   for VITAL
   end for;
end CFG_DLCP1_VITAL;


----- CELL DLCP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := -1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := -1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCP3_3B : entity is TRUE;
end DLCP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLCP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DLCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Tviol_SN_GN_posedge or Pviol_RN or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLCP1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLCP1_QN_tab,
        DataIn => (
               SN_ipd, GN_ipd, RN_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 3 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 3 => (SN_ipd'last_event, tpd_SN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLCP3_VITAL of DLCP3_3B is
   for VITAL
   end for;
end CFG_DLCP3_VITAL;


----- CELL DLCPQ1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCPQ1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCPQ1_3B : entity is TRUE;
end DLCPQ1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLCPQ1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DLCPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Tviol_SN_GN_posedge or Pviol_RN or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLCP1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 3 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLCPQ1_VITAL of DLCPQ1_3B is
   for VITAL
   end for;
end CFG_DLCPQ1_VITAL;


----- CELL DLCPQ3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCPQ3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCPQ3_3B : entity is TRUE;
end DLCPQ3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLCPQ3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/DLCPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Tviol_SN_GN_posedge or Pviol_RN or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLCP1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 3 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLCPQ3_VITAL of DLCPQ3_3B is
   for VITAL
   end for;
end CFG_DLCPQ3_VITAL;


----- CELL DLCQ1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCQ1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCQ1_3B : entity is TRUE;
end DLCQ1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLCQ1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLCQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Pviol_GN or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLCQ1_VITAL of DLCQ1_3B is
   for VITAL
   end for;
end CFG_DLCQ1_VITAL;


----- CELL DLCQ3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCQ3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_RN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCQ3_3B : entity is TRUE;
end DLCQ3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLCQ3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_RN_GN_posedge,
          TimingData              => Tmkr_RN_GN_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_RN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_RN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLCQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_RN_GN_posedge or Pviol_GN or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1_Q_tab,
        DataIn => (
               RN_ipd, GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (RN_ipd'last_event, tpd_RN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLCQ3_VITAL of DLCQ3_3B is
   for VITAL
   end for;
end CFG_DLCQ3_VITAL;


----- CELL DLP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1_3B : entity is TRUE;
end DLP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_SN_GN_posedge or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE),
                 2 => (SN_ipd'last_event, tpd_SN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLP1_VITAL of DLP1_3B is
   for VITAL
   end for;
end CFG_DLP1_VITAL;


----- CELL DLP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := -1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP3_3B : entity is TRUE;
end DLP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_SN_GN_posedge or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_QN, TRUE),
                 2 => (SN_ipd'last_event, tpd_SN_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLP3_VITAL of DLP3_3B is
   for VITAL
   end for;
end CFG_DLP3_VITAL;


----- CELL DLPQ1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLPQ1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLPQ1_3B : entity is TRUE;
end DLPQ1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLPQ1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLPQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_SN_GN_posedge or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLPQ1_VITAL of DLPQ1_3B is
   for VITAL
   end for;
end CFG_DLPQ1_VITAL;


----- CELL DLPQ3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLPQ3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SN_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_GN_posedge_posedge :	VitalDelayType := 0 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of DLPQ3_3B : entity is TRUE;
end DLPQ3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLPQ3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SN_GN_posedge,
          TimingData              => Tmkr_SN_GN_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => trecovery_SN_GN_posedge_posedge,
          SetupLow                => 0 ps,
          HoldHigh                => thold_SN_GN_posedge_posedge,
          HoldLow                 => 0 ps,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLPQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Tviol_SN_GN_posedge or Pviol_GN or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd, SN_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE),
                 2 => (SN_ipd'last_event, tpd_SN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLPQ3_VITAL of DLPQ3_3B is
   for VITAL
   end for;
end CFG_DLPQ3_VITAL;


----- CELL DLQ1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLQ1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLQ1_3B : entity is TRUE;
end DLQ1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLQ1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLQ1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Pviol_GN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLQ1_VITAL of DLQ1_3B is
   for VITAL
   end for;
end CFG_DLQ1_VITAL;


----- CELL DLQ3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLQ3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_GN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_D_GN_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_D_GN_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_D_GN_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_D_GN_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_GN_negedge                 :	VitalDelayType := 1 ps;
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_GN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      D                              :	in    STD_ULOGIC;
      GN                             :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLQ3_3B : entity is TRUE;
end DLQ3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLQ3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (GN_ipd, GN, tipd_GN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, GN_ipd)

   -- timing check results
   VARIABLE Tviol_D_GN_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GN_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GN_posedge,
          TimingData              => Tmkr_D_GN_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ps,
          RefSignal               => GN_ipd,
          RefSignalName          => "GN",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_D_GN_posedge_posedge,
          SetupLow                => tsetup_D_GN_negedge_posedge,
          HoldHigh                => thold_D_GN_posedge_posedge,
          HoldLow                 => thold_D_GN_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GN,
          PeriodData              => PInfo_GN,
          TestSignal              => GN_ipd,
          TestSignalName          => "GN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_GN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLQ3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GN_posedge or Pviol_GN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1_Q_tab,
        DataIn => (
               GN_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (GN_ipd'last_event, tpd_GN_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLQ3_VITAL of DLQ3_3B is
   for VITAL
   end for;
end CFG_DLQ3_VITAL;


----- CELL DLY12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLY12_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLY12_3B : entity is TRUE;
end DLY12_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLY12_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLY12_VITAL of DLY12_3B is
   for VITAL
   end for;
end CFG_DLY12_VITAL;


----- CELL DLY22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLY22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLY22_3B : entity is TRUE;
end DLY22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLY22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLY22_VITAL of DLY22_3B is
   for VITAL
   end for;
end CFG_DLY22_VITAL;


----- CELL DLY32 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLY32_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLY32_3B : entity is TRUE;
end DLY32_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLY32_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLY32_VITAL of DLY32_3B is
   for VITAL
   end for;
end CFG_DLY32_VITAL;


----- CELL DLY42 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLY42_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLY42_3B : entity is TRUE;
end DLY42_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of DLY42_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLY42_VITAL of DLY42_3B is
   for VITAL
   end for;
end CFG_DLY42_VITAL;


----- CELL IMAJ30 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMAJ30_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IMAJ30_3B : entity is TRUE;
end IMAJ30_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMAJ30_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd :=
       (NOT (((B_ipd) AND (C_ipd)) OR ((A_ipd) AND (B_ipd)) OR ((A_ipd) AND
         (C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMAJ30_VITAL of IMAJ30_3B is
   for VITAL
   end for;
end CFG_IMAJ30_VITAL;


----- CELL IMAJ31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMAJ31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IMAJ31_3B : entity is TRUE;
end IMAJ31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMAJ31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd :=
       (NOT (((B_ipd) AND (C_ipd)) OR ((A_ipd) AND (B_ipd)) OR ((A_ipd) AND
         (C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMAJ31_VITAL of IMAJ31_3B is
   for VITAL
   end for;
end CFG_IMAJ31_VITAL;


----- CELL IMUX20 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX20_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX20_3B : entity is TRUE;
end IMUX20_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX20_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX20_VITAL of IMUX20_3B is
   for VITAL
   end for;
end CFG_IMUX20_VITAL;


----- CELL IMUX21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX21_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX21_3B : entity is TRUE;
end IMUX21_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX21_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX21_VITAL of IMUX21_3B is
   for VITAL
   end for;
end CFG_IMUX21_VITAL;


----- CELL IMUX22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX22_3B : entity is TRUE;
end IMUX22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX22_VITAL of IMUX22_3B is
   for VITAL
   end for;
end CFG_IMUX22_VITAL;


----- CELL IMUX23 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX23_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX23_3B : entity is TRUE;
end IMUX23_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX23_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX23_VITAL of IMUX23_3B is
   for VITAL
   end for;
end CFG_IMUX23_VITAL;


----- CELL IMUX24 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX24_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX24_3B : entity is TRUE;
end IMUX24_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX24_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX24_VITAL of IMUX24_3B is
   for VITAL
   end for;
end CFG_IMUX24_VITAL;


----- CELL IMUX30 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX30_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX30_3B : entity is TRUE;
end IMUX30_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX30_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 4 => (S1_ipd'last_event, tpd_S1_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX30_VITAL of IMUX30_3B is
   for VITAL
   end for;
end CFG_IMUX30_VITAL;


----- CELL IMUX31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX31_3B : entity is TRUE;
end IMUX31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 4 => (S1_ipd'last_event, tpd_S1_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX31_VITAL of IMUX31_3B is
   for VITAL
   end for;
end CFG_IMUX31_VITAL;


----- CELL IMUX32 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX32_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX32_3B : entity is TRUE;
end IMUX32_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX32_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 4 => (S1_ipd'last_event, tpd_S1_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX32_VITAL of IMUX32_3B is
   for VITAL
   end for;
end CFG_IMUX32_VITAL;


----- CELL IMUX33 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX33_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX33_3B : entity is TRUE;
end IMUX33_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX33_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 4 => (S1_ipd'last_event, tpd_S1_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX33_VITAL of IMUX33_3B is
   for VITAL
   end for;
end CFG_IMUX33_VITAL;


----- CELL IMUX40 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX40_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX40_3B : entity is TRUE;
end IMUX40_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX40_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (D_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX40_VITAL of IMUX40_3B is
   for VITAL
   end for;
end CFG_IMUX40_VITAL;


----- CELL IMUX41 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX41_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX41_3B : entity is TRUE;
end IMUX41_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX41_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (D_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX41_VITAL of IMUX41_3B is
   for VITAL
   end for;
end CFG_IMUX41_VITAL;


----- CELL IMUX42 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IMUX42_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of IMUX42_3B : entity is TRUE;
end IMUX42_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of IMUX42_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (D_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));
      Q_zd := NOT Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_IMUX42_VITAL of IMUX42_3B is
   for VITAL
   end for;
end CFG_IMUX42_VITAL;


----- CELL INV0 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV0_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV0_3B : entity is TRUE;
end INV0_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV0_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV0_VITAL of INV0_3B is
   for VITAL
   end for;
end CFG_INV0_VITAL;


----- CELL INV1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV1_3B : entity is TRUE;
end INV1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV1_VITAL of INV1_3B is
   for VITAL
   end for;
end CFG_INV1_VITAL;


----- CELL INV2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV2_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV2_3B : entity is TRUE;
end INV2_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV2_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV2_VITAL of INV2_3B is
   for VITAL
   end for;
end CFG_INV2_VITAL;


----- CELL INV3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV3_3B : entity is TRUE;
end INV3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV3_VITAL of INV3_3B is
   for VITAL
   end for;
end CFG_INV3_VITAL;


----- CELL INV4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV4_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV4_3B : entity is TRUE;
end INV4_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV4_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV4_VITAL of INV4_3B is
   for VITAL
   end for;
end CFG_INV4_VITAL;


----- CELL INV6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV6_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV6_3B : entity is TRUE;
end INV6_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV6_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV6_VITAL of INV6_3B is
   for VITAL
   end for;
end CFG_INV6_VITAL;


----- CELL INV8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV8_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV8_3B : entity is TRUE;
end INV8_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV8_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV8_VITAL of INV8_3B is
   for VITAL
   end for;
end CFG_INV8_VITAL;


----- CELL INV10 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV10_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV10_3B : entity is TRUE;
end INV10_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV10_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV10_VITAL of INV10_3B is
   for VITAL
   end for;
end CFG_INV10_VITAL;


----- CELL INV12 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV12_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV12_3B : entity is TRUE;
end INV12_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV12_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV12_VITAL of INV12_3B is
   for VITAL
   end for;
end CFG_INV12_VITAL;


----- CELL INV15 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV15_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV15_3B : entity is TRUE;
end INV15_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of INV15_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_INV15_VITAL of INV15_3B is
   for VITAL
   end for;
end CFG_INV15_VITAL;


----- CELL JK1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JK1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JK1_3B : entity is TRUE;
end JK1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JK1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JK1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JK1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JK1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JK1_Q_tab,
        DataIn => (
               C_delayed, J_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JK1_VITAL of JK1_3B is
   for VITAL
   end for;
end CFG_JK1_VITAL;


----- CELL JK3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JK3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JK3_3B : entity is TRUE;
end JK3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JK3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JK3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JK3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JK3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JK1_Q_tab,
        DataIn => (
               C_delayed, J_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JK3_VITAL of JK3_3B is
   for VITAL
   end for;
end CFG_JK3_VITAL;


----- CELL JKC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKC1_3B : entity is TRUE;
end JKC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, J_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKC1_VITAL of JKC1_3B is
   for VITAL
   end for;
end CFG_JKC1_VITAL;


----- CELL JKC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKC3_3B : entity is TRUE;
end JKC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, J_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKC3_VITAL of JKC3_3B is
   for VITAL
   end for;
end CFG_JKC3_VITAL;


----- CELL JKCP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKCP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKCP1_3B : entity is TRUE;
end JKCP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKCP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/JKCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => JKCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, K_delayed, Q_zd, J_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, J_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKCP1_VITAL of JKCP1_3B is
   for VITAL
   end for;
end CFG_JKCP1_VITAL;


----- CELL JKCP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKCP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKCP3_3B : entity is TRUE;
end JKCP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKCP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/JKCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => JKCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, K_delayed, Q_zd, J_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, J_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKCP3_VITAL of JKCP3_3B is
   for VITAL
   end for;
end CFG_JKCP3_VITAL;


----- CELL JKP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKP1_3B : entity is TRUE;
end JKP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKP1_Q_tab,
        DataIn => (
               C_delayed, J_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKP1_VITAL of JKP1_3B is
   for VITAL
   end for;
end CFG_JKP1_VITAL;


----- CELL JKP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKP3_3B : entity is TRUE;
end JKP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKP1_Q_tab,
        DataIn => (
               C_delayed, J_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKP3_VITAL of JKP3_3B is
   for VITAL
   end for;
end CFG_JKP3_VITAL;


----- CELL JKS1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKS1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := -1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKS1_3B : entity is TRUE;
end JKS1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKS1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKS1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKS1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKS1_VITAL of JKS1_3B is
   for VITAL
   end for;
end CFG_JKS1_VITAL;


----- CELL JKS3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKS3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := -1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKS3_3B : entity is TRUE;
end JKS3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKS3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SE_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKS3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKS1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKS3_VITAL of JKS3_3B is
   for VITAL
   end for;
end CFG_JKS3_VITAL;


----- CELL JKSC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKSC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := -1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKSC1_3B : entity is TRUE;
end JKSC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKSC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKSC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKSC1_VITAL of JKSC1_3B is
   for VITAL
   end for;
end CFG_JKSC1_VITAL;


----- CELL JKSC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKSC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKSC3_3B : entity is TRUE;
end JKSC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKSC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Pviol_C;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKSC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKSC3_VITAL of JKSC3_3B is
   for VITAL
   end for;
end CFG_JKSC3_VITAL;


----- CELL JKSCP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKSCP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKSCP1_3B : entity is TRUE;
end JKSCP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKSCP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => JKSCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, K_delayed, SE_delayed, Q_zd, J_delayed, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKSCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKSCP1_VITAL of JKSCP1_3B is
   for VITAL
   end for;
end CFG_JKSCP1_VITAL;


----- CELL JKSCP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKSCP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKSCP3_3B : entity is TRUE;
end JKSCP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKSCP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_RN_C_posedge or Pviol_RN or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => JKSCP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, K_delayed, SE_delayed, Q_zd, J_delayed, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKSCP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKSCP3_VITAL of JKSCP3_3B is
   for VITAL
   end for;
end CFG_JKSCP3_VITAL;


----- CELL JKSP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKSP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := -1 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKSP1_3B : entity is TRUE;
end JKSP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKSP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKSP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKSP1_VITAL of JKSP1_3B is
   for VITAL
   end for;
end CFG_JKSP1_VITAL;


----- CELL JKSP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKSP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_J_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_J_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_J_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_J_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_K_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_K_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_K_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_K_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_J                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_K                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of JKSP3_3B : entity is TRUE;
end JKSP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of JKSP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, J_ipd, K_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_J_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_C_posedge,
          TimingData              => Tmkr_J_C_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_J_C_posedge_posedge,
          SetupLow                => tsetup_J_C_negedge_posedge,
          HoldHigh                => thold_J_C_posedge_posedge,
          HoldLow                 => thold_J_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_C_posedge,
          TimingData              => Tmkr_K_C_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_K_C_posedge_posedge,
          SetupLow                => tsetup_K_C_negedge_posedge,
          HoldHigh                => thold_K_C_posedge_posedge,
          HoldLow                 => thold_K_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_C_posedge or Tviol_K_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKSP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, J_delayed, SE_delayed, Q_zd, K_delayed, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_JKSP3_VITAL of JKSP3_3B is
   for VITAL
   end for;
end CFG_JKSP3_VITAL;


----- CELL MAJ31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MAJ31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MAJ31_3B : entity is TRUE;
end MAJ31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MAJ31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd :=
       ((B_ipd) AND (C_ipd)) OR ((A_ipd) AND (B_ipd)) OR ((A_ipd) AND
         (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MAJ31_VITAL of MAJ31_3B is
   for VITAL
   end for;
end CFG_MAJ31_VITAL;


----- CELL MAJ32 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MAJ32_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MAJ32_3B : entity is TRUE;
end MAJ32_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MAJ32_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd :=
       ((B_ipd) AND (C_ipd)) OR ((A_ipd) AND (B_ipd)) OR ((A_ipd) AND
         (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MAJ32_VITAL of MAJ32_3B is
   for VITAL
   end for;
end CFG_MAJ32_VITAL;


----- CELL MUX21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX21_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX21_3B : entity is TRUE;
end MUX21_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX21_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX21_VITAL of MUX21_3B is
   for VITAL
   end for;
end CFG_MUX21_VITAL;


----- CELL MUX22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX22_3B : entity is TRUE;
end MUX22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX22_VITAL of MUX22_3B is
   for VITAL
   end for;
end CFG_MUX22_VITAL;


----- CELL MUX24 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX24_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX24_3B : entity is TRUE;
end MUX24_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX24_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX24_VITAL of MUX24_3B is
   for VITAL
   end for;
end CFG_MUX24_VITAL;


----- CELL MUX26 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX26_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX26_3B : entity is TRUE;
end MUX26_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX26_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX26_VITAL of MUX26_3B is
   for VITAL
   end for;
end CFG_MUX26_VITAL;


----- CELL MUX31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX31_3B : entity is TRUE;
end MUX31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 1 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX31_VITAL of MUX31_3B is
   for VITAL
   end for;
end CFG_MUX31_VITAL;


----- CELL MUX32 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX32_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX32_3B : entity is TRUE;
end MUX32_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX32_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 1 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX32_VITAL of MUX32_3B is
   for VITAL
   end for;
end CFG_MUX32_VITAL;


----- CELL MUX33 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX33_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX33_3B : entity is TRUE;
end MUX33_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX33_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 1 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX33_VITAL of MUX33_3B is
   for VITAL
   end for;
end CFG_MUX33_VITAL;


----- CELL MUX34 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX34_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX34_3B : entity is TRUE;
end MUX34_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX34_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (C_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 1 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX34_VITAL of MUX34_3B is
   for VITAL
   end for;
end CFG_MUX34_VITAL;


----- CELL MUX41 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX41_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX41_3B : entity is TRUE;
end MUX41_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX41_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (D_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 1 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 5 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX41_VITAL of MUX41_3B is
   for VITAL
   end for;
end CFG_MUX41_VITAL;


----- CELL MUX42 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX42_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX42_3B : entity is TRUE;
end MUX42_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX42_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (D_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 1 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 5 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX42_VITAL of MUX42_3B is
   for VITAL
   end for;
end CFG_MUX42_VITAL;


----- CELL MUX43 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MUX43_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_S0_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_S1_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S0                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_S1                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of MUX43_3B : entity is TRUE;
end MUX43_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of MUX43_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := VitalMUX
                 (data => (D_ipd, C_ipd, B_ipd, A_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 1 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 5 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_MUX43_VITAL of MUX43_3B is
   for VITAL
   end for;
end CFG_MUX43_VITAL;


----- CELL NAND20 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND20_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND20_3B : entity is TRUE;
end NAND20_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND20_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) AND (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND20_VITAL of NAND20_3B is
   for VITAL
   end for;
end CFG_NAND20_VITAL;


----- CELL NAND21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND21_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND21_3B : entity is TRUE;
end NAND21_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND21_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) AND (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND21_VITAL of NAND21_3B is
   for VITAL
   end for;
end CFG_NAND21_VITAL;


----- CELL NAND22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND22_3B : entity is TRUE;
end NAND22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) AND (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND22_VITAL of NAND22_3B is
   for VITAL
   end for;
end CFG_NAND22_VITAL;


----- CELL NAND23 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND23_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND23_3B : entity is TRUE;
end NAND23_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND23_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) AND (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND23_VITAL of NAND23_3B is
   for VITAL
   end for;
end CFG_NAND23_VITAL;


----- CELL NAND24 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND24_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND24_3B : entity is TRUE;
end NAND24_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND24_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) AND (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND24_VITAL of NAND24_3B is
   for VITAL
   end for;
end CFG_NAND24_VITAL;


----- CELL NAND26 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND26_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND26_3B : entity is TRUE;
end NAND26_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND26_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) AND (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND26_VITAL of NAND26_3B is
   for VITAL
   end for;
end CFG_NAND26_VITAL;


----- CELL NAND28 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND28_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND28_3B : entity is TRUE;
end NAND28_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND28_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) AND (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND28_VITAL of NAND28_3B is
   for VITAL
   end for;
end CFG_NAND28_VITAL;


----- CELL NAND30 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND30_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND30_3B : entity is TRUE;
end NAND30_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND30_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) AND (C_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND30_VITAL of NAND30_3B is
   for VITAL
   end for;
end CFG_NAND30_VITAL;


----- CELL NAND31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND31_3B : entity is TRUE;
end NAND31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) AND (C_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND31_VITAL of NAND31_3B is
   for VITAL
   end for;
end CFG_NAND31_VITAL;


----- CELL NAND32 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND32_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND32_3B : entity is TRUE;
end NAND32_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND32_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) AND (C_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND32_VITAL of NAND32_3B is
   for VITAL
   end for;
end CFG_NAND32_VITAL;


----- CELL NAND33 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND33_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND33_3B : entity is TRUE;
end NAND33_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND33_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) AND (C_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND33_VITAL of NAND33_3B is
   for VITAL
   end for;
end CFG_NAND33_VITAL;


----- CELL NAND34 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND34_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND34_3B : entity is TRUE;
end NAND34_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND34_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) AND (C_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND34_VITAL of NAND34_3B is
   for VITAL
   end for;
end CFG_NAND34_VITAL;


----- CELL NAND40 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND40_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND40_3B : entity is TRUE;
end NAND40_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND40_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) AND (D_ipd) AND (B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND40_VITAL of NAND40_3B is
   for VITAL
   end for;
end CFG_NAND40_VITAL;


----- CELL NAND41 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND41_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND41_3B : entity is TRUE;
end NAND41_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND41_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) AND (D_ipd) AND (B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND41_VITAL of NAND41_3B is
   for VITAL
   end for;
end CFG_NAND41_VITAL;


----- CELL NAND42 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND42_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND42_3B : entity is TRUE;
end NAND42_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND42_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) AND (D_ipd) AND (B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND42_VITAL of NAND42_3B is
   for VITAL
   end for;
end CFG_NAND42_VITAL;


----- CELL NAND43 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND43_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND43_3B : entity is TRUE;
end NAND43_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NAND43_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) AND (D_ipd) AND (B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NAND43_VITAL of NAND43_3B is
   for VITAL
   end for;
end CFG_NAND43_VITAL;


----- CELL NOR20 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR20_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR20_3B : entity is TRUE;
end NOR20_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR20_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) OR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR20_VITAL of NOR20_3B is
   for VITAL
   end for;
end CFG_NOR20_VITAL;


----- CELL NOR21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR21_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR21_3B : entity is TRUE;
end NOR21_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR21_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) OR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR21_VITAL of NOR21_3B is
   for VITAL
   end for;
end CFG_NOR21_VITAL;


----- CELL NOR22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR22_3B : entity is TRUE;
end NOR22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) OR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR22_VITAL of NOR22_3B is
   for VITAL
   end for;
end CFG_NOR22_VITAL;


----- CELL NOR23 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR23_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR23_3B : entity is TRUE;
end NOR23_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR23_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) OR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR23_VITAL of NOR23_3B is
   for VITAL
   end for;
end CFG_NOR23_VITAL;


----- CELL NOR24 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR24_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR24_3B : entity is TRUE;
end NOR24_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR24_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) OR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR24_VITAL of NOR24_3B is
   for VITAL
   end for;
end CFG_NOR24_VITAL;


----- CELL NOR30 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR30_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR30_3B : entity is TRUE;
end NOR30_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR30_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) OR (C_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR30_VITAL of NOR30_3B is
   for VITAL
   end for;
end CFG_NOR30_VITAL;


----- CELL NOR31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR31_3B : entity is TRUE;
end NOR31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) OR (C_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR31_VITAL of NOR31_3B is
   for VITAL
   end for;
end CFG_NOR31_VITAL;


----- CELL NOR32 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR32_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR32_3B : entity is TRUE;
end NOR32_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR32_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) OR (C_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR32_VITAL of NOR32_3B is
   for VITAL
   end for;
end CFG_NOR32_VITAL;


----- CELL NOR33 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR33_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR33_3B : entity is TRUE;
end NOR33_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR33_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) OR (C_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR33_VITAL of NOR33_3B is
   for VITAL
   end for;
end CFG_NOR33_VITAL;


----- CELL NOR40 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR40_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR40_3B : entity is TRUE;
end NOR40_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR40_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR (D_ipd) OR (B_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR40_VITAL of NOR40_3B is
   for VITAL
   end for;
end CFG_NOR40_VITAL;


----- CELL NOR41 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR41_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR41_3B : entity is TRUE;
end NOR41_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR41_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR (D_ipd) OR (B_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR41_VITAL of NOR41_3B is
   for VITAL
   end for;
end CFG_NOR41_VITAL;


----- CELL NOR42 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR42_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR42_3B : entity is TRUE;
end NOR42_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of NOR42_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) OR (D_ipd) OR (B_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_NOR42_VITAL of NOR42_3B is
   for VITAL
   end for;
end CFG_NOR42_VITAL;


----- CELL OAI210 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI210_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI210_3B : entity is TRUE;
end OAI210_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI210_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((B_ipd) OR (A_ipd)) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI210_VITAL of OAI210_3B is
   for VITAL
   end for;
end CFG_OAI210_VITAL;


----- CELL OAI211 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI211_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI211_3B : entity is TRUE;
end OAI211_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI211_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((B_ipd) OR (A_ipd)) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI211_VITAL of OAI211_3B is
   for VITAL
   end for;
end CFG_OAI211_VITAL;


----- CELL OAI212 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI212_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI212_3B : entity is TRUE;
end OAI212_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI212_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((B_ipd) OR (A_ipd)) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI212_VITAL of OAI212_3B is
   for VITAL
   end for;
end CFG_OAI212_VITAL;


----- CELL OAI220 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI220_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI220_3B : entity is TRUE;
end OAI220_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI220_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((A_ipd) OR (B_ipd)) AND ((C_ipd) OR (D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI220_VITAL of OAI220_3B is
   for VITAL
   end for;
end CFG_OAI220_VITAL;


----- CELL OAI221 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI221_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI221_3B : entity is TRUE;
end OAI221_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI221_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((A_ipd) OR (B_ipd)) AND ((C_ipd) OR (D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI221_VITAL of OAI221_3B is
   for VITAL
   end for;
end CFG_OAI221_VITAL;


----- CELL OAI222 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI222_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI222_3B : entity is TRUE;
end OAI222_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI222_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((A_ipd) OR (B_ipd)) AND ((C_ipd) OR (D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI222_VITAL of OAI222_3B is
   for VITAL
   end for;
end CFG_OAI222_VITAL;


----- CELL OAI310 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI310_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI310_3B : entity is TRUE;
end OAI310_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI310_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((A_ipd) OR (B_ipd) OR (C_ipd)) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI310_VITAL of OAI310_3B is
   for VITAL
   end for;
end CFG_OAI310_VITAL;


----- CELL OAI311 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI311_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI311_3B : entity is TRUE;
end OAI311_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI311_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((A_ipd) OR (B_ipd) OR (C_ipd)) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI311_VITAL of OAI311_3B is
   for VITAL
   end for;
end CFG_OAI311_VITAL;


----- CELL OAI312 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI312_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI312_3B : entity is TRUE;
end OAI312_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI312_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT (((A_ipd) OR (B_ipd) OR (C_ipd)) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI312_VITAL of OAI312_3B is
   for VITAL
   end for;
end CFG_OAI312_VITAL;


----- CELL OAI2110 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI2110_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI2110_3B : entity is TRUE;
end OAI2110_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI2110_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) AND (D_ipd) AND ((A_ipd) OR (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI2110_VITAL of OAI2110_3B is
   for VITAL
   end for;
end CFG_OAI2110_VITAL;


----- CELL OAI2111 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI2111_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI2111_3B : entity is TRUE;
end OAI2111_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI2111_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) AND (D_ipd) AND ((A_ipd) OR (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI2111_VITAL of OAI2111_3B is
   for VITAL
   end for;
end CFG_OAI2111_VITAL;


----- CELL OAI2112 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI2112_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI2112_3B : entity is TRUE;
end OAI2112_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of OAI2112_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) AND (D_ipd) AND ((A_ipd) OR (B_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_OAI2112_VITAL of OAI2112_3B is
   for VITAL
   end for;
end CFG_OAI2112_VITAL;


----- CELL TFC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFC1_3B : entity is TRUE;
end TFC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFC1_VITAL of TFC1_3B is
   for VITAL
   end for;
end CFG_TFC1_VITAL;


----- CELL TFC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFC3_3B : entity is TRUE;
end TFC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFC3_VITAL of TFC3_3B is
   for VITAL
   end for;
end CFG_TFC3_VITAL;


----- CELL TFCP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFCP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFCP1_3B : entity is TRUE;
end TFCP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFCP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFCP1_Q_tab,
        DataIn => (
               SN_ipd, C_delayed, Q_zd, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFCP1_QN_tab,
        DataIn => (
               RN_ipd, C_delayed, SN_ipd, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFCP1_VITAL of TFCP1_3B is
   for VITAL
   end for;
end CFG_TFCP1_VITAL;


----- CELL TFCP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFCP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFCP3_3B : entity is TRUE;
end TFCP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFCP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFCP1_Q_tab,
        DataIn => (
               SN_ipd, C_delayed, Q_zd, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFCP1_QN_tab,
        DataIn => (
               RN_ipd, C_delayed, SN_ipd, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFCP3_VITAL of TFCP3_3B is
   for VITAL
   end for;
end CFG_TFCP3_VITAL;


----- CELL TFEC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFEC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFEC1_3B : entity is TRUE;
end TFEC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFEC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_T_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, T_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFEC1_VITAL of TFEC1_3B is
   for VITAL
   end for;
end CFG_TFEC1_VITAL;


----- CELL TFEC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFEC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFEC3_3B : entity is TRUE;
end TFEC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFEC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_T_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, T_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFEC3_VITAL of TFEC3_3B is
   for VITAL
   end for;
end CFG_TFEC3_VITAL;


----- CELL TFECP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFECP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFECP1_3B : entity is TRUE;
end TFECP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFECP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => TFECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, T_delayed, Q_zd, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFECP1_VITAL of TFECP1_3B is
   for VITAL
   end for;
end CFG_TFECP1_VITAL;


----- CELL TFECP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFECP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFECP3_3B : entity is TRUE;
end TFECP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFECP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => TFECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, T_delayed, Q_zd, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFECP3_VITAL of TFECP3_3B is
   for VITAL
   end for;
end CFG_TFECP3_VITAL;


----- CELL TFEP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFEP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFEP1_3B : entity is TRUE;
end TFEP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFEP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SN_C_posedge or Pviol_C or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFEP1_Q_tab,
        DataIn => (
               C_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFEP1_VITAL of TFEP1_3B is
   for VITAL
   end for;
end CFG_TFEP1_VITAL;


----- CELL TFEP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFEP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := -1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFEP3_3B : entity is TRUE;
end TFEP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFEP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SN_C_posedge or Pviol_C or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFEP1_Q_tab,
        DataIn => (
               C_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFEP3_VITAL of TFEP3_3B is
   for VITAL
   end for;
end CFG_TFEP3_VITAL;


----- CELL TFP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFP1_3B : entity is TRUE;
end TFP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFP1_Q_tab,
        DataIn => (
               C_delayed, SN_ipd, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFP1_VITAL of TFP1_3B is
   for VITAL
   end for;
end CFG_TFP1_VITAL;


----- CELL TFP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFP3_3B : entity is TRUE;
end TFP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFP1_Q_tab,
        DataIn => (
               C_delayed, SN_ipd, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFP3_VITAL of TFP3_3B is
   for VITAL
   end for;
end CFG_TFP3_VITAL;


----- CELL TFSC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSC1_3B : entity is TRUE;
end TFSC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSC1_VITAL of TFSC1_3B is
   for VITAL
   end for;
end CFG_TFSC1_VITAL;


----- CELL TFSC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSC3_3B : entity is TRUE;
end TFSC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSC3_VITAL of TFSC3_3B is
   for VITAL
   end for;
end CFG_TFSC3_VITAL;


----- CELL TFSCP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSCP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSCP1_3B : entity is TRUE;
end TFSCP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSCP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSCP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => JKCP1_Q_tab,
        DataIn => (
               SN_ipd, C_delayed, Q_zd, SE_delayed, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKCP1_QN_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSCP1_VITAL of TFSCP1_3B is
   for VITAL
   end for;
end CFG_TFSCP1_VITAL;


----- CELL TFSCP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSCP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSCP3_3B : entity is TRUE;
end TFSCP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSCP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSCP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => JKCP1_Q_tab,
        DataIn => (
               SN_ipd, C_delayed, Q_zd, SE_delayed, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => JKCP1_QN_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSCP3_VITAL of TFSCP3_3B is
   for VITAL
   end for;
end CFG_TFSCP3_VITAL;


----- CELL TFSEC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSEC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := -1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSEC1_3B : entity is TRUE;
end TFSEC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSEC1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSEC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_T_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, T_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSEC1_VITAL of TFSEC1_3B is
   for VITAL
   end for;
end CFG_TFSEC1_VITAL;


----- CELL TFSEC3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSEC3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_RN_Q                       :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := 1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := -1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSEC3_3B : entity is TRUE;
end TFSEC3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSEC3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT RN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSEC3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_T_C_posedge or Pviol_C or Pviol_RN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSEC1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, T_delayed, Q_zd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_RN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSEC3_VITAL of TFSEC3_3B is
   for VITAL
   end for;
end CFG_TFSEC3_VITAL;


----- CELL TFSECP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSECP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSECP1_3B : entity is TRUE;
end TFSECP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSECP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSECP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => TFSECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, SE_delayed, T_delayed, Q_zd, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSECP1_VITAL of TFSECP1_3B is
   for VITAL
   end for;
end CFG_TFSECP1_VITAL;


----- CELL TFSECP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSECP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_RN_Q                       :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_RN_QN                      :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      trecovery_RN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_RN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_RN_negedge                 :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_RN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      RN                             :	in    STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSECP3_3B : entity is TRUE;
end TFSECP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSECP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL RN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (RN_ipd, RN, tipd_RN);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, RN_ipd, SD_ipd, SE_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_RN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_RN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_RN	: STD_ULOGIC := '0';
   VARIABLE PInfo_RN	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_RN_C_posedge,
          TimingData              => Tmkr_RN_C_posedge,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_RN_C_posedge_posedge,
          Removal                 => thold_RN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR ( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT SN_ipd) ) OR ( (NOT RN_ipd) ) ) /=
                            '1',
          HeaderMsg               => InstancePath &"/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_RN,
          PeriodData              => PInfo_RN,
          TestSignal              => RN_ipd,
          TestSignalName          => "RN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_RN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSECP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_RN_C_posedge or Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_RN or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => TFSECP1_QN_tab,
        DataIn => (
               SN_ipd, C_delayed, SE_delayed, T_delayed, Q_zd, SD_delayed, RN_ipd, C_ipd));
      QN_zd := Violation XOR QN_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSECP1_Q_tab,
        DataIn => (
               RN_ipd, C_delayed, SD_delayed, SE_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (RN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (SN_ipd'last_event, tpd_RN_QN, TRUE),
                 2 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSECP3_VITAL of TFSECP3_3B is
   for VITAL
   end for;
end CFG_TFSECP3_VITAL;


----- CELL TFSEP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSEP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSEP1_3B : entity is TRUE;
end TFSEP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSEP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SD_ipd, SE_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSEP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSEP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, SE_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSEP1_VITAL of TFSEP1_3B is
   for VITAL
   end for;
end CFG_TFSEP1_VITAL;


----- CELL TFSEP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSEP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := -1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_T_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_T_C_negedge_posedge      :	VitalDelayType := 1 ps;
      tsetup_T_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_T_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_T                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC;
      T                              :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSEP3_3B : entity is TRUE;
end TFSEP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSEP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL T_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   VitalWireDelay (T_ipd, T, tipd_T);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SD_ipd, SE_ipd, SN_ipd, T_ipd)

   -- timing check results
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_T_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_T_C_posedge,
          TimingData              => Tmkr_T_C_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_T_C_posedge_posedge,
          SetupLow                => tsetup_T_C_negedge_posedge,
          HoldHigh                => thold_T_C_posedge_posedge,
          HoldLow                 => thold_T_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSEP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Tviol_T_C_posedge or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSEP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, SE_delayed, T_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;
      T_delayed := T_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSEP3_VITAL of TFSEP3_3B is
   for VITAL
   end for;
end CFG_TFSEP3_VITAL;


----- CELL TFSP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSP1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSP1_3B : entity is TRUE;
end TFSP1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSP1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, SE_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSP1_VITAL of TFSP1_3B is
   for VITAL
   end for;
end CFG_TFSP1_VITAL;


----- CELL TFSP3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TFSP3_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_SN_Q                       :	VitalDelayType01 := (1 ps, 0 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_SN_QN                      :	VitalDelayType01 := (0 ps, 1 ps);
      tpd_C_QN                       :	VitalDelayType01 := (1 ps, 1 ps);
      thold_SD_C_posedge_posedge     :	VitalDelayType := -1 ps;
      thold_SD_C_negedge_posedge     :	VitalDelayType := -1 ps;
      tsetup_SD_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SD_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := -1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 0 ps;
      trecovery_SN_C_posedge_posedge :	VitalDelayType := 0 ps;
      thold_SN_C_posedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_posedge                  :	VitalDelayType := 1 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tpw_SN_negedge                 :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SD                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SN                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC;
      QN                             :	out   STD_ULOGIC;
      SD                             :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      SN                             :	in    STD_ULOGIC);
attribute VITAL_LEVEL0 of TFSP3_3B : entity is TRUE;
end TFSP3_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TFSP3_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (SD_ipd, SD, tipd_SD);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   VitalWireDelay (SN_ipd, SN, tipd_SN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, SD_ipd, SE_ipd, SN_ipd)

   -- timing check results
   VARIABLE Tviol_SD_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SD_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SN_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SN_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_SN	: STD_ULOGIC := '0';
   VARIABLE PInfo_SN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE C_delayed : STD_ULOGIC := 'X';
   VARIABLE SD_delayed : STD_ULOGIC := 'X';
   VARIABLE SE_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);
   ALIAS QN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_SD_C_posedge,
          TimingData              => Tmkr_SD_C_posedge,
          TestSignal              => SD_ipd,
          TestSignalName          => "SD",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SD_C_posedge_posedge,
          SetupLow                => tsetup_SD_C_negedge_posedge,
          HoldHigh                => thold_SD_C_posedge_posedge,
          HoldLow                 => thold_SD_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT SE_ipd) OR (NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_SN_C_posedge,
          TimingData              => Tmkr_SN_C_posedge,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          Recovery                => trecovery_SN_C_posedge_posedge,
          Removal                 => thold_SN_C_posedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => tpw_C_posedge,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TO_X01((NOT SN_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_SN,
          PeriodData              => PInfo_SN,
          TestSignal              => SN_ipd,
          TestSignalName          => "SN",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_SN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TFSP3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_SD_C_posedge or Tviol_SE_C_posedge or Tviol_SN_C_posedge or Pviol_C or Pviol_SN;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TFSP1_Q_tab,
        DataIn => (
               C_delayed, SD_delayed, SE_delayed, Q_zd, SN_ipd, C_ipd));
      Q_zd := Violation XOR Q_zd;
      QN_zd := (NOT Q_zd);
      C_delayed := C_ipd;
      SD_delayed := SD_ipd;
      SE_delayed := SE_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_Q, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (SN_ipd'last_event, tpd_SN_QN, TRUE),
                 1 => (C_ipd'last_event, tpd_C_QN, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_TFSP3_VITAL of TFSP3_3B is
   for VITAL
   end for;
end CFG_TFSP3_VITAL;


----- CELL TIE0 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TIE0_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True);

   port(
      Q                              :	out   STD_ULOGIC := '0');
attribute VITAL_LEVEL0 of TIE0_3B : entity is TRUE;
end TIE0_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TIE0_3B is
   attribute VITAL_LEVEL0 of VITAL : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Q <= '0';


end VITAL;

configuration CFG_TIE0_VITAL of TIE0_3B is
   for VITAL
   end for;
end CFG_TIE0_VITAL;


----- CELL TIE1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TIE1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True);

   port(
      Q                              :	out   STD_ULOGIC := '1');
attribute VITAL_LEVEL0 of TIE1_3B : entity is TRUE;
end TIE1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of TIE1_3B is
   attribute VITAL_LEVEL0 of VITAL : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Q <= '1';


end VITAL;

configuration CFG_TIE1_VITAL of TIE1_3B is
   for VITAL
   end for;
end CFG_TIE1_VITAL;


----- CELL XNR20 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNR20_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNR20_3B : entity is TRUE;
end XNR20_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XNR20_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) XOR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XNR20_VITAL of XNR20_3B is
   for VITAL
   end for;
end CFG_XNR20_VITAL;


----- CELL XNR21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNR21_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNR21_3B : entity is TRUE;
end XNR21_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XNR21_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) XOR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XNR21_VITAL of XNR21_3B is
   for VITAL
   end for;
end CFG_XNR21_VITAL;


----- CELL XNR22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNR22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNR22_3B : entity is TRUE;
end XNR22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XNR22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((A_ipd) XOR (B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XNR22_VITAL of XNR22_3B is
   for VITAL
   end for;
end CFG_XNR22_VITAL;


----- CELL XNR30 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNR30_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNR30_3B : entity is TRUE;
end XNR30_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XNR30_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) XOR (C_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XNR30_VITAL of XNR30_3B is
   for VITAL
   end for;
end CFG_XNR30_VITAL;


----- CELL XNR31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNR31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNR31_3B : entity is TRUE;
end XNR31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XNR31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((B_ipd) XOR (C_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XNR31_VITAL of XNR31_3B is
   for VITAL
   end for;
end CFG_XNR31_VITAL;


----- CELL XNR40 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNR40_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNR40_3B : entity is TRUE;
end XNR40_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XNR40_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) XOR (D_ipd) XOR (B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XNR40_VITAL of XNR40_3B is
   for VITAL
   end for;
end CFG_XNR40_VITAL;


----- CELL XNR41 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNR41_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNR41_3B : entity is TRUE;
end XNR41_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XNR41_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (NOT ((C_ipd) XOR (D_ipd) XOR (B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XNR41_VITAL of XNR41_3B is
   for VITAL
   end for;
end CFG_XNR41_VITAL;


----- CELL XOR20 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR20_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR20_3B : entity is TRUE;
end XOR20_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XOR20_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (A_ipd) XOR (B_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XOR20_VITAL of XOR20_3B is
   for VITAL
   end for;
end CFG_XOR20_VITAL;


----- CELL XOR21 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR21_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR21_3B : entity is TRUE;
end XOR21_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XOR21_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (A_ipd) XOR (B_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XOR21_VITAL of XOR21_3B is
   for VITAL
   end for;
end CFG_XOR21_VITAL;


----- CELL XOR22 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR22_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR22_3B : entity is TRUE;
end XOR22_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XOR22_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (A_ipd) XOR (B_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XOR22_VITAL of XOR22_3B is
   for VITAL
   end for;
end CFG_XOR22_VITAL;


----- CELL XOR30 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR30_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR30_3B : entity is TRUE;
end XOR30_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XOR30_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (B_ipd) XOR (C_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XOR30_VITAL of XOR30_3B is
   for VITAL
   end for;
end CFG_XOR30_VITAL;


----- CELL XOR31 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR31_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR31_3B : entity is TRUE;
end XOR31_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XOR31_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (B_ipd) XOR (C_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XOR31_VITAL of XOR31_3B is
   for VITAL
   end for;
end CFG_XOR31_VITAL;


----- CELL XOR40 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR40_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR40_3B : entity is TRUE;
end XOR40_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XOR40_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (C_ipd) XOR (D_ipd) XOR (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XOR40_VITAL of XOR40_3B is
   for VITAL
   end for;
end CFG_XOR40_VITAL;


----- CELL XOR41 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR41_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_B_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_C_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tpd_D_Q                        :	VitalDelayType01 := (1 ps, 1 ps);
      tipd_A                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_B                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_D                         :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR41_3B : entity is TRUE;
end XOR41_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB_3B;
use c35_CORELIB_3B.VTABLES.all;
architecture VITAL of XOR41_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Q_zd := (C_ipd) XOR (D_ipd) XOR (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Q, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Q, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_XOR41_VITAL of XOR41_3B is
   for VITAL
   end for;
end CFG_XOR41_VITAL;


----- CELL DLSG1_3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLSG1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_C_GCK                      :	VitalDelayType01 := (1 ps, 1 ps);
      tsetup_E_C_posedge_posedge     :	VitalDelayType := 1 ps;
      tsetup_E_C_negedge_posedge     :	VitalDelayType := 1 ps;
      thold_E_C_posedge_posedge      :	VitalDelayType := 0 ps;
      thold_E_C_negedge_posedge      :	VitalDelayType := 0 ps;
      tsetup_SE_C_posedge_posedge    :	VitalDelayType := 1 ps;
      tsetup_SE_C_negedge_posedge    :	VitalDelayType := 1 ps;
      thold_SE_C_posedge_posedge     :	VitalDelayType := 0 ps;
      thold_SE_C_negedge_posedge     :	VitalDelayType := 0 ps;
      tpw_C_negedge                  :	VitalDelayType := 1 ps;
      tipd_C                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_E                         :	VitalDelayType01 := (0 ps, 0 ps);
      tipd_SE                        :	VitalDelayType01 := (0 ps, 0 ps));

   port(
      C                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      SE                             :	in    STD_ULOGIC;
      GCK                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLSG1_3B : entity is TRUE;
end DLSG1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB;
use c35_CORELIB.VTABLES.all;
architecture VITAL of DLSG1_3B is
   attribute VITAL_LEVEL1 of VITAL : architecture is TRUE;

   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL SE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (SE_ipd, SE, tipd_SE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (C_ipd, E_ipd, SE_ipd)

   -- timing check results
   VARIABLE Tviol_E_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_SE_C_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_SE_C_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_C	: STD_ULOGIC := '0';
   VARIABLE PInfo_C	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_IQ : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE IQ : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS GCK_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE GCK_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_E_C_posedge,
          TimingData              => Tmkr_E_C_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_E_C_posedge_posedge,
          SetupLow                => tsetup_E_C_negedge_posedge,
          HoldHigh                => thold_E_C_posedge_posedge,
          HoldLow                 => thold_E_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLSG1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_SE_C_posedge,
          TimingData              => Tmkr_SE_C_posedge,
          TestSignal              => SE_ipd,
          TestSignalName          => "SE",
          TestDelay               => 0 ps,
          RefSignal               => C_ipd,
          RefSignalName          => "C",
          RefDelay                => 0 ps,
          SetupHigh               => tsetup_SE_C_posedge_posedge,
          SetupLow                => tsetup_SE_C_negedge_posedge,
          HoldHigh                => thold_SE_C_posedge_posedge,
          HoldLow                 => thold_SE_C_negedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLSG1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_C,
          PeriodData              => PInfo_C,
          TestSignal              => C_ipd,
          TestSignalName          => "C",
          TestDelay               => 0 ps,
          Period                  => 0 ps,
          PulseWidthHigh          => 0 ps,
          PulseWidthLow           => tpw_C_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLSG1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_E_C_posedge or Pviol_C or Tviol_SE_C_posedge;
      VitalStateTable(
        Result => IQ,
        PreviousDataIn => PrevData_IQ,
        StateTable => DLSG1_IQ_tab,
        DataIn => (
               C_ipd, SE_ipd, E_ipd));
      IQ := Violation XOR IQ;
      GCK_zd := (C_ipd) AND (IQ);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => GCK,
       GlitchData => GCK_GlitchData,
       OutSignalName => "GCK",
       OutTemp => GCK_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_GCK, TRUE)),
       Mode => OnEvent,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL;

configuration CFG_DLSG1_VITAL of DLSG1_3B is
   for VITAL
   end for;
end CFG_DLSG1_VITAL;


----- CELL LOGIC0_3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity LOGIC0_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True);

   port(
      Q                              :	out   STD_ULOGIC := '0');
attribute VITAL_LEVEL0 of LOGIC0_3B : entity is TRUE;
end LOGIC0_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB;
use c35_CORELIB.VTABLES.all;
architecture VITAL of LOGIC0_3B is
   attribute VITAL_LEVEL0 of VITAL : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Q <= '0';


end VITAL;

configuration CFG_LOGIC0_VITAL of LOGIC0_3B is
   for VITAL
   end for;
end CFG_LOGIC0_VITAL;


----- CELL LOGIC1_3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity LOGIC1_3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True);

   port(
      Q                              :	out   STD_ULOGIC := '1');
attribute VITAL_LEVEL0 of LOGIC1_3B : entity is TRUE;
end LOGIC1_3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library c35_CORELIB;
use c35_CORELIB.VTABLES.all;
architecture VITAL of LOGIC1_3B is
   attribute VITAL_LEVEL0 of VITAL : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Q <= '1';


end VITAL;

configuration CFG_LOGIC1_VITAL of LOGIC1_3B is
   for VITAL
   end for;
end CFG_LOGIC1_VITAL;




---- end of library ----

