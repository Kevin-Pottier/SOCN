library IEEE;
use IEEE.electrical_systems.all;
use IEEE.math_real.all;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity bod_vhdlams is
  port(terminal tvdd,tvss,tbod_det,tbod_en : ELECTRICAL);
  end entity bod_vhdlams;

library ieee;
use ieee.math_real.all;

architecture behav of bod_vhdlams is
begin

end architecture behav;

