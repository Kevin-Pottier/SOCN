//-------------------------------------------------------------------------
// ﾩ 1997-2005 Cadence Design Systems, Inc.  All rights reserved.
// This work may not be copied, modified, re-published, uploaded, executed,
// or distributed in any way, in any medium, whether in whole or in part,
// without prior written permission from Cadence Design Systems, Inc.
//------------------------------------------------------------------------

//------------------------------------------------------------------------
//  Abstract   : Simulation Architecture for v06
//  RC Release : v06.20-s026_1
//------------------------------------------------------------------------


module GTECH_FD2S (D, CP, TI, TE, CD, Q, QN);  
	input D, CP, CD, TI, TE;
	output Q, QN;

	reg Q, QN;
	
	always @(Q)
        begin
                QN = ~Q;
        end

        always @(posedge CP or negedge CD)
        begin
	    begin
	    	if (!CD)
		    Q = 1'b0;
	        else if (TE)
		    Q = TI;
	    	else
                    Q = D;
	    end
        end
endmodule



